library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


entity rom is
	port(
		clock:   in  std_logic;
		rd_addr: in  std_logic_vector(7 downto 0);
		q:       out std_logic_vector(7 downto 0)
	);
end rom;


architecture a of rom is
	type mem is array(0 to 255) of std_logic_vector(7 downto 0);
	signal storage: mem := (
		b"00001000", 
		b"00001000", 
		b"00010000", 
		b"00001000", 
		b"00010000", 
		b"00001000", 
		b"00000100", 
		b"00000100", 
		b"00001000", 
		b"00010000", 
		b"00100000", 
		b"00100000", 
		b"00010000", 
		b"00001000", 
		b"00000100", 
		b"00000010", 
		b"00000010", 
		b"00000100", 
		b"00001000", 
		b"00010000", 
		b"00100000", 
		b"01000000", 
		b"01000000", 
		b"00100000", 
		b"00010000", 
		b"00001000", 
		b"00000100", 
		b"00000010", 
		b"00000001", 
		b"00000001", 
		b"00000010", 
		b"00000100", 
		b"00001000", 
		b"00010000", 
		b"00100000", 
		b"01000000", 
		b"10000000", 
		b"10000000", 
		b"10000000", 
		b"01000000", 
		b"00100000", 
		b"00010000", 
		b"00001000", 
		b"00000100", 
		b"00000010", 
		b"00000010", 
		b"00000010", 
		b"00000101", 
		b"00001000", 
		b"00001000", 
		b"00010000", 
		b"00001000", 
		b"00010000", 
		b"00001000", 
		b"00000100", 
		b"00000100", 
		b"00001000", 
		b"00010000", 
		b"00100000", 
		b"00100000", 
		b"00010000", 
		b"00001000", 
		b"00000100", 
		b"00000010", 
		b"00000010", 
		b"00000100", 
		b"00001000", 
		b"00010000", 
		b"00100000", 
		b"01000000", 
		b"01000000", 
		b"00100000", 
		b"00010000", 
		b"00001000", 
		b"00000100", 
		b"00000010", 
		b"00000001", 
		b"00000001", 
		b"00000010", 
		b"00000100", 
		b"00001000", 
		b"00010000", 
		b"00100000", 
		b"01000000", 
		b"10000000", 
		b"10000000", 
		b"10000000", 
		b"01000000", 
		b"00100000", 
		b"00010000", 
		b"00001000", 
		b"00000100", 
		b"00000010", 
		b"00000001", 
		b"00000001", 
		b"00000001", 
		b"00001000", 
		b"00001000", 
		b"00010000", 
		b"00001000", 
		b"00010000", 
		b"00001000", 
		b"00000100", 
		b"00000100", 
		b"00001000", 
		b"00010000", 
		b"00100000", 
		b"00100000", 
		b"00010000", 
		b"00001000", 
		b"00000100", 
		b"00000010", 
		b"00000010", 
		b"00000100", 
		b"00001000", 
		b"00010000", 
		b"00100000", 
		b"01000000", 
		b"01000000", 
		b"00100000", 
		b"00010000", 
		b"00001000", 
		b"00000100", 
		b"00000010", 
		b"00000001", 
		b"00000001", 
		b"00000010", 
		b"00000100", 
		b"00001000", 
		b"00010000", 
		b"00100000", 
		b"01000000", 
		b"10000000", 
		b"10000000", 
		b"10000000", 
		b"01000000", 
		b"00100000", 
		b"00010000", 
		b"00001000", 
		b"00000100", 
		b"00000010", 
		b"00000010", 
		b"00000010", 
		b"00000101", 
		b"00001000", 
		b"00001000", 
		b"00010000", 
		b"00001000", 
		b"00010000", 
		b"00001000", 
		b"00000100", 
		b"00000100", 
		b"00001000", 
		b"00010000", 
		b"00100000", 
		b"00100000", 
		b"00010000", 
		b"00001000", 
		b"00000100", 
		b"00000010", 
		b"00000010", 
		b"00000100", 
		b"00001000", 
		b"00010000", 
		b"00100000", 
		b"01000000", 
		b"01000000", 
		b"00100000", 
		b"00010000", 
		b"00001000", 
		b"00000100", 
		b"00000010", 
		b"00000001", 
		b"00000001", 
		b"00000010", 
		b"00000100", 
		b"00001000", 
		b"00010000", 
		b"00100000", 
		b"01000000", 
		b"10000000", 
		b"10000000", 
		b"10000000", 
		b"01000000", 
		b"00100000", 
		b"00010000", 
		b"00001000", 
		b"00000100", 
		b"00000010", 
		b"00000001", 
		b"00000001", 
		b"00000001",
		b"00000010", 
		b"00000010", 
		b"00000100", 
		b"00001000", 
		b"00010000", 
		b"00100000", 
		b"01000000", 
		b"01000000", 
		b"00100000", 
		b"00010000", 
		b"00001000", 
		b"00000100", 
		b"00000010", 
		b"00000001", 
		b"00000001", 
		b"00000010", 
		b"00000100", 
		b"00001000", 
		b"00010000", 
		b"00100000", 
		b"01000000", 
		b"10000000", 
		b"10000000", 
		b"10000000", 
		b"01000000", 
		b"00100000", 
		b"00010000", 
		b"00001000", 
		b"00000100", 
		b"00000010", 
		b"00000001", 
		b"00000010", 
		b"00000100",
		b"00001000",
		b"00001000", 
		b"00010000", 
		b"00100000", 
		b"01000000", 
		b"01000000", 
		b"00100000", 
		b"00010000", 
		b"00001000", 
		b"00000100", 
		b"00000010", 
		b"00000001", 
		b"00000001", 
		b"00000010", 
		b"00000100", 
		b"00001000", 
		b"00010000", 
		b"00100000", 
		b"01000000", 
		b"10000000", 
		b"10000000", 
		b"10000000", 
		b"01000000", 
		b"00100000", 
		b"00010000", 
		b"00001000", 
		b"00000100", 
		b"00000010", 
		b"00000001", 
		b"00000010", 
		b"00001000"
	);
begin

	q <= storage(to_integer(unsigned(rd_addr))) when rising_edge(clock);

end a;
